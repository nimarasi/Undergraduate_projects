library verilog;
use verilog.vl_types.all;
entity FullAdder_vlg_vec_tst is
end FullAdder_vlg_vec_tst;
