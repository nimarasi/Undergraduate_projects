library verilog;
use verilog.vl_types.all;
entity full_vlg_vec_tst is
end full_vlg_vec_tst;
