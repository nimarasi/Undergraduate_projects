library verilog;
use verilog.vl_types.all;
entity b2g_vlg_vec_tst is
end b2g_vlg_vec_tst;
