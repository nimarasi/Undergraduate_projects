library verilog;
use verilog.vl_types.all;
entity encoder_vlg_check_tst is
    port(
        y0              : in     vl_logic;
        y1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end encoder_vlg_check_tst;
