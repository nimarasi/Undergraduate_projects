library verilog;
use verilog.vl_types.all;
entity bu_vlg_vec_tst is
end bu_vlg_vec_tst;
